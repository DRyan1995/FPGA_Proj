`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:02:37 12/22/2015 
// Design Name: 
// Module Name:    sigtap 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sigtap( touch_in,touch_out
    );
	 input touch_in;
	 output touch_out;
	 assign touch_out=touch_in;


endmodule
