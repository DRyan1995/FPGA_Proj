`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:15:04 12/23/2015 
// Design Name: 
// Module Name:    MP3 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MP3(
		inout mp3_in,
		inout mp3_out
    );
	
	assign mp3_out = mp3_in;
		

endmodule
