// CORE V2.v

// Generated using ACDS version 13.0 156 at 2015.12.19.13:37:15

`timescale 1 ps / 1 ps
module CORE V2 (
		input  wire        clk_clk,                        //                       clk.clk
		input  wire        reset_reset_n,                  //                     reset.reset_n
		input  wire        rs232_external_connection_rxd,  // rs232_external_connection.rxd
		output wire        rs232_external_connection_txd,  //                          .txd
		output wire [11:0] sdram_controller_wire_addr,     //     sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,       //                          .ba
		output wire        sdram_controller_wire_cas_n,    //                          .cas_n
		output wire        sdram_controller_wire_cke,      //                          .cke
		output wire        sdram_controller_wire_cs_n,     //                          .cs_n
		inout  wire [15:0] sdram_controller_wire_dq,       //                          .dq
		output wire [1:0]  sdram_controller_wire_dqm,      //                          .dqm
		output wire        sdram_controller_wire_ras_n,    //                          .ras_n
		output wire        sdram_controller_wire_we_n,     //                          .we_n
		output wire [7:0]  out_external_connection_export, //   out_external_connection.export
		input  wire [3:0]  in_external_connection_export   //    in_external_connection.export
	);

	wire         nios2_instruction_master_waitrequest;                                                             // nios2_instruction_master_translator:av_waitrequest -> nios2:i_waitrequest
	wire  [24:0] nios2_instruction_master_address;                                                                 // nios2:i_address -> nios2_instruction_master_translator:av_address
	wire         nios2_instruction_master_read;                                                                    // nios2:i_read -> nios2_instruction_master_translator:av_read
	wire  [31:0] nios2_instruction_master_readdata;                                                                // nios2_instruction_master_translator:av_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_readdatavalid;                                                           // nios2_instruction_master_translator:av_readdatavalid -> nios2:i_readdatavalid
	wire         nios2_data_master_waitrequest;                                                                    // nios2_data_master_translator:av_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                                                                      // nios2:d_writedata -> nios2_data_master_translator:av_writedata
	wire  [24:0] nios2_data_master_address;                                                                        // nios2:d_address -> nios2_data_master_translator:av_address
	wire         nios2_data_master_write;                                                                          // nios2:d_write -> nios2_data_master_translator:av_write
	wire         nios2_data_master_read;                                                                           // nios2:d_read -> nios2_data_master_translator:av_read
	wire  [31:0] nios2_data_master_readdata;                                                                       // nios2_data_master_translator:av_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                                                                    // nios2:jtag_debug_module_debugaccess_to_roms -> nios2_data_master_translator:av_debugaccess
	wire         nios2_data_master_readdatavalid;                                                                  // nios2_data_master_translator:av_readdatavalid -> nios2:d_readdatavalid
	wire   [3:0] nios2_data_master_byteenable;                                                                     // nios2:d_byteenable -> nios2_data_master_translator:av_byteenable
	wire         nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                               // nios2:jtag_debug_module_waitrequest -> nios2_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                 // nios2_jtag_debug_module_translator:av_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_address;                                   // nios2_jtag_debug_module_translator:av_address -> nios2:jtag_debug_module_address
	wire         nios2_jtag_debug_module_translator_avalon_anti_slave_0_write;                                     // nios2_jtag_debug_module_translator:av_write -> nios2:jtag_debug_module_write
	wire         nios2_jtag_debug_module_translator_avalon_anti_slave_0_read;                                      // nios2_jtag_debug_module_translator:av_read -> nios2:jtag_debug_module_read
	wire  [31:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                  // nios2:jtag_debug_module_readdata -> nios2_jtag_debug_module_translator:av_readdata
	wire         nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                               // nios2_jtag_debug_module_translator:av_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                // nios2_jtag_debug_module_translator:av_byteenable -> nios2:jtag_debug_module_byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire   [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire         sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest;                                   // sdram_controller:za_waitrequest -> sdram_controller_s1_translator:av_waitrequest
	wire  [15:0] sdram_controller_s1_translator_avalon_anti_slave_0_writedata;                                     // sdram_controller_s1_translator:av_writedata -> sdram_controller:az_data
	wire  [21:0] sdram_controller_s1_translator_avalon_anti_slave_0_address;                                       // sdram_controller_s1_translator:av_address -> sdram_controller:az_addr
	wire         sdram_controller_s1_translator_avalon_anti_slave_0_chipselect;                                    // sdram_controller_s1_translator:av_chipselect -> sdram_controller:az_cs
	wire         sdram_controller_s1_translator_avalon_anti_slave_0_write;                                         // sdram_controller_s1_translator:av_write -> sdram_controller:az_wr_n
	wire         sdram_controller_s1_translator_avalon_anti_slave_0_read;                                          // sdram_controller_s1_translator:av_read -> sdram_controller:az_rd_n
	wire  [15:0] sdram_controller_s1_translator_avalon_anti_slave_0_readdata;                                      // sdram_controller:za_data -> sdram_controller_s1_translator:av_readdata
	wire         sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid;                                 // sdram_controller:za_valid -> sdram_controller_s1_translator:av_readdatavalid
	wire   [1:0] sdram_controller_s1_translator_avalon_anti_slave_0_byteenable;                                    // sdram_controller_s1_translator:av_byteenable -> sdram_controller:az_be_n
	wire   [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                       // sysid_control_slave_translator:av_address -> sysid:address
	wire  [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                      // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire  [15:0] rs232_s1_translator_avalon_anti_slave_0_writedata;                                                // RS232_s1_translator:av_writedata -> RS232:writedata
	wire   [2:0] rs232_s1_translator_avalon_anti_slave_0_address;                                                  // RS232_s1_translator:av_address -> RS232:address
	wire         rs232_s1_translator_avalon_anti_slave_0_chipselect;                                               // RS232_s1_translator:av_chipselect -> RS232:chipselect
	wire         rs232_s1_translator_avalon_anti_slave_0_write;                                                    // RS232_s1_translator:av_write -> RS232:write_n
	wire         rs232_s1_translator_avalon_anti_slave_0_read;                                                     // RS232_s1_translator:av_read -> RS232:read_n
	wire  [15:0] rs232_s1_translator_avalon_anti_slave_0_readdata;                                                 // RS232:readdata -> RS232_s1_translator:av_readdata
	wire         rs232_s1_translator_avalon_anti_slave_0_begintransfer;                                            // RS232_s1_translator:av_begintransfer -> RS232:begintransfer
	wire  [31:0] myout_s1_translator_avalon_anti_slave_0_writedata;                                                // MYOUT_s1_translator:av_writedata -> MYOUT:writedata
	wire   [1:0] myout_s1_translator_avalon_anti_slave_0_address;                                                  // MYOUT_s1_translator:av_address -> MYOUT:address
	wire         myout_s1_translator_avalon_anti_slave_0_chipselect;                                               // MYOUT_s1_translator:av_chipselect -> MYOUT:chipselect
	wire         myout_s1_translator_avalon_anti_slave_0_write;                                                    // MYOUT_s1_translator:av_write -> MYOUT:write_n
	wire  [31:0] myout_s1_translator_avalon_anti_slave_0_readdata;                                                 // MYOUT:readdata -> MYOUT_s1_translator:av_readdata
	wire   [1:0] myin_s1_translator_avalon_anti_slave_0_address;                                                   // MYIN_s1_translator:av_address -> MYIN:address
	wire  [31:0] myin_s1_translator_avalon_anti_slave_0_readdata;                                                  // MYIN:readdata -> MYIN_s1_translator:av_readdata
	wire         nios2_instruction_master_translator_avalon_universal_master_0_waitrequest;                        // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_instruction_master_translator_avalon_universal_master_0_burstcount;                         // nios2_instruction_master_translator:uav_burstcount -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_instruction_master_translator_avalon_universal_master_0_writedata;                          // nios2_instruction_master_translator:uav_writedata -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] nios2_instruction_master_translator_avalon_universal_master_0_address;                            // nios2_instruction_master_translator:uav_address -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_instruction_master_translator_avalon_universal_master_0_lock;                               // nios2_instruction_master_translator:uav_lock -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_instruction_master_translator_avalon_universal_master_0_write;                              // nios2_instruction_master_translator:uav_write -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_instruction_master_translator_avalon_universal_master_0_read;                               // nios2_instruction_master_translator:uav_read -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_instruction_master_translator_avalon_universal_master_0_readdata;                           // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_instruction_master_translator:uav_readdata
	wire         nios2_instruction_master_translator_avalon_universal_master_0_debugaccess;                        // nios2_instruction_master_translator:uav_debugaccess -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_instruction_master_translator_avalon_universal_master_0_byteenable;                         // nios2_instruction_master_translator:uav_byteenable -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid;                      // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_instruction_master_translator:uav_readdatavalid
	wire         nios2_data_master_translator_avalon_universal_master_0_waitrequest;                               // nios2_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_data_master_translator_avalon_universal_master_0_burstcount;                                // nios2_data_master_translator:uav_burstcount -> nios2_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_data_master_translator_avalon_universal_master_0_writedata;                                 // nios2_data_master_translator:uav_writedata -> nios2_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] nios2_data_master_translator_avalon_universal_master_0_address;                                   // nios2_data_master_translator:uav_address -> nios2_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_data_master_translator_avalon_universal_master_0_lock;                                      // nios2_data_master_translator:uav_lock -> nios2_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_data_master_translator_avalon_universal_master_0_write;                                     // nios2_data_master_translator:uav_write -> nios2_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_data_master_translator_avalon_universal_master_0_read;                                      // nios2_data_master_translator:uav_read -> nios2_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_data_master_translator_avalon_universal_master_0_readdata;                                  // nios2_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_data_master_translator:uav_readdata
	wire         nios2_data_master_translator_avalon_universal_master_0_debugaccess;                               // nios2_data_master_translator:uav_debugaccess -> nios2_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_data_master_translator_avalon_universal_master_0_byteenable;                                // nios2_data_master_translator:uav_byteenable -> nios2_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_data_master_translator_avalon_universal_master_0_readdatavalid;                             // nios2_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_data_master_translator:uav_readdatavalid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // nios2_jtag_debug_module_translator:uav_waitrequest -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                   // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_jtag_debug_module_translator:uav_writedata
	wire  [24:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                     // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_jtag_debug_module_translator:uav_address
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                       // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_jtag_debug_module_translator:uav_write
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                        // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_jtag_debug_module_translator:uav_lock
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                        // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                    // nios2_jtag_debug_module_translator:uav_readdata -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // nios2_jtag_debug_module_translator:uav_readdatavalid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_jtag_debug_module_translator:uav_byteenable
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                 // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire  [24:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // sdram_controller_s1_translator:uav_waitrequest -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_controller_s1_translator:uav_burstcount
	wire  [15:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_controller_s1_translator:uav_writedata
	wire  [24:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_controller_s1_translator:uav_address
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_controller_s1_translator:uav_write
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_controller_s1_translator:uav_lock
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_controller_s1_translator:uav_read
	wire  [15:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // sdram_controller_s1_translator:uav_readdata -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // sdram_controller_s1_translator:uav_readdatavalid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_controller_s1_translator:uav_debugaccess
	wire   [1:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_controller_s1_translator:uav_byteenable
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [80:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [80:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [17:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;               // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [17:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;               // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire  [24:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // RS232_s1_translator:uav_waitrequest -> RS232_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // RS232_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> RS232_s1_translator:uav_burstcount
	wire  [31:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // RS232_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> RS232_s1_translator:uav_writedata
	wire  [24:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // RS232_s1_translator_avalon_universal_slave_0_agent:m0_address -> RS232_s1_translator:uav_address
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // RS232_s1_translator_avalon_universal_slave_0_agent:m0_write -> RS232_s1_translator:uav_write
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // RS232_s1_translator_avalon_universal_slave_0_agent:m0_lock -> RS232_s1_translator:uav_lock
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // RS232_s1_translator_avalon_universal_slave_0_agent:m0_read -> RS232_s1_translator:uav_read
	wire  [31:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // RS232_s1_translator:uav_readdata -> RS232_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // RS232_s1_translator:uav_readdatavalid -> RS232_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // RS232_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RS232_s1_translator:uav_debugaccess
	wire   [3:0] rs232_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // RS232_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> RS232_s1_translator:uav_byteenable
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // RS232_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // RS232_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // RS232_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // RS232_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RS232_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RS232_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RS232_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RS232_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RS232_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // RS232_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // RS232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RS232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // RS232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RS232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // RS232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RS232_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         myout_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // MYOUT_s1_translator:uav_waitrequest -> MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] myout_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> MYOUT_s1_translator:uav_burstcount
	wire  [31:0] myout_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> MYOUT_s1_translator:uav_writedata
	wire  [24:0] myout_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_address -> MYOUT_s1_translator:uav_address
	wire         myout_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_write -> MYOUT_s1_translator:uav_write
	wire         myout_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_lock -> MYOUT_s1_translator:uav_lock
	wire         myout_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_read -> MYOUT_s1_translator:uav_read
	wire  [31:0] myout_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // MYOUT_s1_translator:uav_readdata -> MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         myout_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // MYOUT_s1_translator:uav_readdatavalid -> MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         myout_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> MYOUT_s1_translator:uav_debugaccess
	wire   [3:0] myout_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // MYOUT_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> MYOUT_s1_translator:uav_byteenable
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] myout_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // MYOUT_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // MYOUT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> MYOUT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] myout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // MYOUT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> MYOUT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // MYOUT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> MYOUT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         myin_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // MYIN_s1_translator:uav_waitrequest -> MYIN_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] myin_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // MYIN_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> MYIN_s1_translator:uav_burstcount
	wire  [31:0] myin_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // MYIN_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> MYIN_s1_translator:uav_writedata
	wire  [24:0] myin_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // MYIN_s1_translator_avalon_universal_slave_0_agent:m0_address -> MYIN_s1_translator:uav_address
	wire         myin_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // MYIN_s1_translator_avalon_universal_slave_0_agent:m0_write -> MYIN_s1_translator:uav_write
	wire         myin_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // MYIN_s1_translator_avalon_universal_slave_0_agent:m0_lock -> MYIN_s1_translator:uav_lock
	wire         myin_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // MYIN_s1_translator_avalon_universal_slave_0_agent:m0_read -> MYIN_s1_translator:uav_read
	wire  [31:0] myin_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // MYIN_s1_translator:uav_readdata -> MYIN_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         myin_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // MYIN_s1_translator:uav_readdatavalid -> MYIN_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         myin_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // MYIN_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> MYIN_s1_translator:uav_debugaccess
	wire   [3:0] myin_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // MYIN_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> MYIN_s1_translator:uav_byteenable
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // MYIN_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // MYIN_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // MYIN_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] myin_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // MYIN_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> MYIN_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> MYIN_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> MYIN_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> MYIN_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> MYIN_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // MYIN_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // MYIN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> MYIN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] myin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // MYIN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> MYIN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // MYIN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> MYIN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;               // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                     // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;             // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [97:0] nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                      // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router:sink_ready -> nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // nios2_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid;                            // nios2_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // nios2_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [97:0] nios2_data_master_translator_avalon_universal_master_0_agent_cp_data;                             // nios2_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_001:sink_ready -> nios2_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                       // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [97:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                        // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router:sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [97:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_001:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [79:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_002:sink_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [97:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_003:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // RS232_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // RS232_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // RS232_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [97:0] rs232_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // RS232_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         rs232_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_004:sink_ready -> RS232_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // MYOUT_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // MYOUT_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // MYOUT_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [97:0] myout_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // MYOUT_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         myout_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_005:sink_ready -> MYOUT_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // MYIN_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // MYIN_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // MYIN_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [97:0] myin_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // MYIN_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         myin_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_006:sink_ready -> MYIN_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                      // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                            // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                    // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [97:0] addr_router_src_data;                                                                             // addr_router:src_data -> limiter:cmd_sink_data
	wire   [6:0] addr_router_src_channel;                                                                          // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                            // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                      // limiter:rsp_src_endofpacket -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                            // limiter:rsp_src_valid -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                    // limiter:rsp_src_startofpacket -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [97:0] limiter_rsp_src_data;                                                                             // limiter:rsp_src_data -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [6:0] limiter_rsp_src_channel;                                                                          // limiter:rsp_src_channel -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                            // nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                  // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                        // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [97:0] addr_router_001_src_data;                                                                         // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [6:0] addr_router_001_src_channel;                                                                      // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                        // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                  // limiter_001:rsp_src_endofpacket -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                        // limiter_001:rsp_src_valid -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                // limiter_001:rsp_src_startofpacket -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [97:0] limiter_001_rsp_src_data;                                                                         // limiter_001:rsp_src_data -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [6:0] limiter_001_rsp_src_channel;                                                                      // limiter_001:rsp_src_channel -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                        // nios2_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         burst_adapter_source0_endofpacket;                                                                // burst_adapter:source0_endofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                      // burst_adapter:source0_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                              // burst_adapter:source0_startofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [79:0] burst_adapter_source0_data;                                                                       // burst_adapter:source0_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                      // sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [6:0] burst_adapter_source0_channel;                                                                    // burst_adapter:source0_channel -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                   // rst_controller:reset_out -> [MYIN:reset_n, MYIN_s1_translator:reset, MYIN_s1_translator_avalon_universal_slave_0_agent:reset, MYIN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, MYOUT:reset_n, MYOUT_s1_translator:reset, MYOUT_s1_translator_avalon_universal_slave_0_agent:reset, MYOUT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RS232:reset_n, RS232_s1_translator:reset, RS232_s1_translator_avalon_universal_slave_0_agent:reset, RS232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2:reset_n, nios2_data_master_translator:reset, nios2_data_master_translator_avalon_universal_master_0_agent:reset, nios2_instruction_master_translator:reset, nios2_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_jtag_debug_module_translator:reset, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram_controller:reset_n, sdram_controller_s1_translator:reset, sdram_controller_s1_translator_avalon_universal_slave_0_agent:reset, sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire         nios2_jtag_debug_module_reset_reset;                                                              // nios2:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         cmd_xbar_demux_src0_endofpacket;                                                                  // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                        // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src0_data;                                                                         // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [6:0] cmd_xbar_demux_src0_channel;                                                                      // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                        // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                  // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                        // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src1_data;                                                                         // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [6:0] cmd_xbar_demux_src1_channel;                                                                      // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                        // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                  // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                        // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src2_data;                                                                         // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [6:0] cmd_xbar_demux_src2_channel;                                                                      // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                        // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src0_data;                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [6:0] cmd_xbar_demux_001_src0_channel;                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                    // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                              // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                    // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                            // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src1_data;                                                                     // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [6:0] cmd_xbar_demux_001_src1_channel;                                                                  // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                    // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                              // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                    // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                            // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src2_data;                                                                     // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [6:0] cmd_xbar_demux_001_src2_channel;                                                                  // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                    // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                              // cmd_xbar_demux_001:src3_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                    // cmd_xbar_demux_001:src3_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                            // cmd_xbar_demux_001:src3_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src3_data;                                                                     // cmd_xbar_demux_001:src3_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_001_src3_channel;                                                                  // cmd_xbar_demux_001:src3_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                              // cmd_xbar_demux_001:src4_endofpacket -> RS232_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                    // cmd_xbar_demux_001:src4_valid -> RS232_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                            // cmd_xbar_demux_001:src4_startofpacket -> RS232_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src4_data;                                                                     // cmd_xbar_demux_001:src4_data -> RS232_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_001_src4_channel;                                                                  // cmd_xbar_demux_001:src4_channel -> RS232_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                              // cmd_xbar_demux_001:src5_endofpacket -> MYOUT_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                    // cmd_xbar_demux_001:src5_valid -> MYOUT_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                            // cmd_xbar_demux_001:src5_startofpacket -> MYOUT_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src5_data;                                                                     // cmd_xbar_demux_001:src5_data -> MYOUT_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_001_src5_channel;                                                                  // cmd_xbar_demux_001:src5_channel -> MYOUT_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                              // cmd_xbar_demux_001:src6_endofpacket -> MYIN_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                    // cmd_xbar_demux_001:src6_valid -> MYIN_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                            // cmd_xbar_demux_001:src6_startofpacket -> MYIN_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src6_data;                                                                     // cmd_xbar_demux_001:src6_data -> MYIN_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_001_src6_channel;                                                                  // cmd_xbar_demux_001:src6_channel -> MYIN_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                  // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                        // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [97:0] rsp_xbar_demux_src0_data;                                                                         // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [6:0] rsp_xbar_demux_src0_channel;                                                                      // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                        // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                  // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                        // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [97:0] rsp_xbar_demux_src1_data;                                                                         // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [6:0] rsp_xbar_demux_src1_channel;                                                                      // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                        // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                              // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                    // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                            // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [97:0] rsp_xbar_demux_001_src0_data;                                                                     // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [6:0] rsp_xbar_demux_001_src0_channel;                                                                  // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                    // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                              // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                    // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                            // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [97:0] rsp_xbar_demux_001_src1_data;                                                                     // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [6:0] rsp_xbar_demux_001_src1_channel;                                                                  // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                    // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                              // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                    // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                            // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [97:0] rsp_xbar_demux_002_src0_data;                                                                     // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [6:0] rsp_xbar_demux_002_src0_channel;                                                                  // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                    // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                              // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                    // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                            // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [97:0] rsp_xbar_demux_002_src1_data;                                                                     // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [6:0] rsp_xbar_demux_002_src1_channel;                                                                  // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                    // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                              // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                    // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                            // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [97:0] rsp_xbar_demux_003_src0_data;                                                                     // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [6:0] rsp_xbar_demux_003_src0_channel;                                                                  // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                    // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                              // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                    // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                            // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [97:0] rsp_xbar_demux_004_src0_data;                                                                     // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [6:0] rsp_xbar_demux_004_src0_channel;                                                                  // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                    // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                              // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                    // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                            // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [97:0] rsp_xbar_demux_005_src0_data;                                                                     // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [6:0] rsp_xbar_demux_005_src0_channel;                                                                  // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                    // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                              // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                    // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                            // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [97:0] rsp_xbar_demux_006_src0_data;                                                                     // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [6:0] rsp_xbar_demux_006_src0_channel;                                                                  // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                    // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                      // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                    // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [97:0] limiter_cmd_src_data;                                                                             // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [6:0] limiter_cmd_src_channel;                                                                          // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                            // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                     // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                           // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                   // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [97:0] rsp_xbar_mux_src_data;                                                                            // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [6:0] rsp_xbar_mux_src_channel;                                                                         // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                           // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                  // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [97:0] limiter_001_cmd_src_data;                                                                         // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [6:0] limiter_001_cmd_src_channel;                                                                      // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                        // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                 // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                       // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                               // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [97:0] rsp_xbar_mux_001_src_data;                                                                        // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [6:0] rsp_xbar_mux_001_src_channel;                                                                     // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                       // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                     // cmd_xbar_mux:src_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                           // cmd_xbar_mux:src_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                   // cmd_xbar_mux:src_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_src_data;                                                                            // cmd_xbar_mux:src_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_mux_src_channel;                                                                         // cmd_xbar_mux:src_channel -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                           // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [97:0] id_router_src_data;                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [6:0] id_router_src_channel;                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                 // cmd_xbar_mux_001:src_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                       // cmd_xbar_mux_001:src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                               // cmd_xbar_mux_001:src_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_001_src_data;                                                                        // cmd_xbar_mux_001:src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_mux_001_src_channel;                                                                     // cmd_xbar_mux_001:src_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                    // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                          // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                  // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [97:0] id_router_001_src_data;                                                                           // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [6:0] id_router_001_src_channel;                                                                        // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                          // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                    // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                          // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                  // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [97:0] id_router_003_src_data;                                                                           // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [6:0] id_router_003_src_channel;                                                                        // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                          // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                    // RS232_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                    // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                          // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                  // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [97:0] id_router_004_src_data;                                                                           // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [6:0] id_router_004_src_channel;                                                                        // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                          // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                    // MYOUT_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                    // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                          // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                  // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [97:0] id_router_005_src_data;                                                                           // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [6:0] id_router_005_src_channel;                                                                        // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                          // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                    // MYIN_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                    // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                          // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                  // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [97:0] id_router_006_src_data;                                                                           // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [6:0] id_router_006_src_channel;                                                                        // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                          // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                 // cmd_xbar_mux_002:src_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                       // cmd_xbar_mux_002:src_valid -> width_adapter:in_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                               // cmd_xbar_mux_002:src_startofpacket -> width_adapter:in_startofpacket
	wire  [97:0] cmd_xbar_mux_002_src_data;                                                                        // cmd_xbar_mux_002:src_data -> width_adapter:in_data
	wire   [6:0] cmd_xbar_mux_002_src_channel;                                                                     // cmd_xbar_mux_002:src_channel -> width_adapter:in_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                       // width_adapter:in_ready -> cmd_xbar_mux_002:src_ready
	wire         width_adapter_src_endofpacket;                                                                    // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                          // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                  // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [79:0] width_adapter_src_data;                                                                           // width_adapter:out_data -> burst_adapter:sink0_data
	wire         width_adapter_src_ready;                                                                          // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [6:0] width_adapter_src_channel;                                                                        // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire         id_router_002_src_endofpacket;                                                                    // id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_002_src_valid;                                                                          // id_router_002:src_valid -> width_adapter_001:in_valid
	wire         id_router_002_src_startofpacket;                                                                  // id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [79:0] id_router_002_src_data;                                                                           // id_router_002:src_data -> width_adapter_001:in_data
	wire   [6:0] id_router_002_src_channel;                                                                        // id_router_002:src_channel -> width_adapter_001:in_channel
	wire         id_router_002_src_ready;                                                                          // width_adapter_001:in_ready -> id_router_002:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                // width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                      // width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                              // width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [97:0] width_adapter_001_src_data;                                                                       // width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	wire         width_adapter_001_src_ready;                                                                      // rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	wire   [6:0] width_adapter_001_src_channel;                                                                    // width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	wire   [6:0] limiter_cmd_valid_data;                                                                           // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [6:0] limiter_001_cmd_valid_data;                                                                       // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                         // RS232:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                         // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_d_irq_irq;                                                                                  // irq_mapper:sender_irq -> nios2:d_irq

	CORE V2_nios2 nios2 (
		.clk                                   (clk_clk),                                                            //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                    //                   reset_n.reset_n
		.d_address                             (nios2_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_data_master_writedata),                                        //                          .writedata
		.d_readdatavalid                       (nios2_data_master_readdatavalid),                                    //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	CORE V2_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                //               irq.irq
	);

	CORE V2_RS232 rs232 (
		.clk           (clk_clk),                                               //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address       (rs232_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (rs232_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (rs232_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~rs232_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~rs232_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (rs232_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (rs232_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                      //                    .dataavailable
		.readyfordata  (),                                                      //                    .readyfordata
		.rxd           (rs232_external_connection_rxd),                         // external_connection.export
		.txd           (rs232_external_connection_txd),                         //                    .export
		.irq           (irq_mapper_receiver0_irq)                               //                 irq.irq
	);

	CORE V2_sysid sysid (
		.clock    (clk_clk),                                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	CORE V2_sdram_controller sdram_controller (
		.clk            (clk_clk),                                                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                                  // reset.reset_n
		.az_addr        (sdram_controller_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_controller_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_controller_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_controller_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_controller_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_controller_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_controller_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_controller_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_controller_wire_dq),                                         //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                                        //      .export
	);

	CORE V2_MYOUT myout (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (myout_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~myout_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (myout_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (myout_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (myout_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_external_connection_export)                      // external_connection.export
	);

	CORE V2_MYIN myin (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (myin_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (myin_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (in_external_connection_export)                    // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_instruction_master_translator (
		.clk                      (clk_clk),                                                                     //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_byteenable            (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_write                 (1'b0),                                                                        //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_data_master_translator (
		.clk                      (clk_clk),                                                              //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address              (nios2_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_data_master_read),                                               //                          .read
		.av_readdata              (nios2_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (nios2_data_master_write),                                              //                          .write
		.av_writedata             (nios2_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_chipselect            (1'b0),                                                                 //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_chipselect            (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_controller_s1_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_controller_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_controller_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_controller_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_controller_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_controller_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_controller_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_controller_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rs232_s1_translator (
		.clk                      (clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (rs232_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (rs232_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (rs232_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (rs232_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (rs232_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (rs232_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (rs232_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (rs232_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (rs232_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (rs232_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (rs232_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (rs232_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (rs232_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (rs232_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (rs232_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (rs232_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) myout_s1_translator (
		.clk                      (clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (myout_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (myout_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (myout_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (myout_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (myout_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (myout_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (myout_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (myout_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (myout_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (myout_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (myout_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (myout_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (myout_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (myout_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (myout_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (myout_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) myin_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (myin_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (myin_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (myin_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (myin_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (myin_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (myin_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (myin_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (myin_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (myin_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (myin_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (myin_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (myin_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (myin_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                   //              (terminated)
		.av_read                  (),                                                                   //              (terminated)
		.av_writedata             (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_chipselect            (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_THREAD_ID_H           (88),
		.PKT_THREAD_ID_L           (88),
		.PKT_CACHE_H               (95),
		.PKT_CACHE_L               (92),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.ST_DATA_W                 (98),
		.ST_CHANNEL_W              (7),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                              //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                                //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                                 //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                              //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                        //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                          //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                                //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_THREAD_ID_H           (88),
		.PKT_THREAD_ID_L           (88),
		.PKT_CACHE_H               (95),
		.PKT_CACHE_L               (92),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.ST_DATA_W                 (98),
		.ST_CHANNEL_W              (7),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                       //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address              (nios2_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                     //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                      //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                   //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                             //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                               //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                     //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                                     //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (62),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (66),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (67),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_controller_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                              //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                              //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                               //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                        //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                            //                .channel
		.rf_sink_ready           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_startofpacket  (1'b0),                                                                               // (terminated)
		.in_endofpacket    (1'b0),                                                                               // (terminated)
		.out_startofpacket (),                                                                                   // (terminated)
		.out_endofpacket   (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) rs232_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (rs232_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rs232_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rs232_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rs232_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rs232_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rs232_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rs232_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rs232_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rs232_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rs232_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rs232_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rs232_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rs232_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rs232_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rs232_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                               //                .channel
		.rf_sink_ready           (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rs232_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rs232_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rs232_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) myout_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (myout_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (myout_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (myout_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (myout_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (myout_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (myout_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (myout_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (myout_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (myout_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (myout_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (myout_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (myout_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (myout_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (myout_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (myout_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (myout_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                               //                .channel
		.rf_sink_ready           (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (myout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (myout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (myout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (myout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (myout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (myout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (myout_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (myout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) myin_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (myin_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (myin_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (myin_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (myin_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (myin_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (myin_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (myin_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (myin_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (myin_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (myin_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (myin_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (myin_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (myin_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (myin_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (myin_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (myin_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                              //                .channel
		.rf_sink_ready           (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (myin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (myin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (myin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (myin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (myin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (myin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (myin_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (myin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	CORE V2_addr_router addr_router (
		.sink_ready         (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	CORE V2_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	CORE V2_id_router id_router (
		.sink_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	CORE V2_id_router id_router_001 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                //          .valid
		.src_data           (id_router_001_src_data),                                                                 //          .data
		.src_channel        (id_router_001_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                           //          .endofpacket
	);

	CORE V2_id_router_002 id_router_002 (
		.sink_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                        //       src.ready
		.src_valid          (id_router_002_src_valid),                                                        //          .valid
		.src_data           (id_router_002_src_data),                                                         //          .data
		.src_channel        (id_router_002_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                   //          .endofpacket
	);

	CORE V2_id_router_003 id_router_003 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                        //       src.ready
		.src_valid          (id_router_003_src_valid),                                                        //          .valid
		.src_data           (id_router_003_src_data),                                                         //          .data
		.src_channel        (id_router_003_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                   //          .endofpacket
	);

	CORE V2_id_router_003 id_router_004 (
		.sink_ready         (rs232_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rs232_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rs232_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rs232_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rs232_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                             //       src.ready
		.src_valid          (id_router_004_src_valid),                                             //          .valid
		.src_data           (id_router_004_src_data),                                              //          .data
		.src_channel        (id_router_004_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                        //          .endofpacket
	);

	CORE V2_id_router_003 id_router_005 (
		.sink_ready         (myout_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (myout_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (myout_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (myout_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (myout_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                             //       src.ready
		.src_valid          (id_router_005_src_valid),                                             //          .valid
		.src_data           (id_router_005_src_data),                                              //          .data
		.src_channel        (id_router_005_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                        //          .endofpacket
	);

	CORE V2_id_router_003 id_router_006 (
		.sink_ready         (myin_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (myin_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (myin_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (myin_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (myin_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                            //       src.ready
		.src_valid          (id_router_006_src_valid),                                            //          .valid
		.src_data           (id_router_006_src_data),                                             //          .data
		.src_channel        (id_router_006_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                       //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (98),
		.ST_CHANNEL_W              (7),
		.VALID_WIDTH               (7),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (98),
		.ST_CHANNEL_W              (7),
		.VALID_WIDTH               (7),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (62),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.PKT_BURST_TYPE_H          (59),
		.PKT_BURST_TYPE_L          (58),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (7),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (54),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clk_clk),                             //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	CORE V2_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //           .endofpacket
	);

	CORE V2_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket)    //           .endofpacket
	);

	CORE V2_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	CORE V2_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	CORE V2_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	CORE V2_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	CORE V2_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	CORE V2_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	CORE V2_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	CORE V2_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	CORE V2_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	CORE V2_rsp_xbar_demux_003 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	CORE V2_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	CORE V2_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (69),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (70),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (97),
		.IN_PKT_RESPONSE_STATUS_L      (96),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (98),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (51),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (57),
		.OUT_PKT_BURST_SIZE_L          (55),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (59),
		.OUT_PKT_BURST_TYPE_L          (58),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clk_clk),                            //       clk.clk
		.reset                (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_mux_002_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_002_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_002_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_002_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_002_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (51),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (54),
		.IN_PKT_BURSTWRAP_L            (52),
		.IN_PKT_BURST_SIZE_H           (57),
		.IN_PKT_BURST_SIZE_L           (55),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (59),
		.IN_PKT_BURST_TYPE_L           (58),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (69),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (97),
		.OUT_PKT_RESPONSE_STATUS_L     (96),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (98),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_002_src_valid),             //      sink.valid
		.in_channel           (id_router_002_src_channel),           //          .channel
		.in_startofpacket     (id_router_002_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_002_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_002_src_ready),             //          .ready
		.in_data              (id_router_002_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	CORE V2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

endmodule
